`define ADDR_WIDTH 8
`define DATA_WIDTH 16
`define DEPTH 256
`define RESET_VAL 16'h1234

import uvm_pkg::*;