class test extends uvm_test;
    `uvm_component_utils(test)
    function new(string name = "test", uvm_component parent=null);
      super.new(name, parent);
    endfunction
  
    env e0;
    virtual reg_if vif;

    // virtual function void start_of_simulation_phase(uvm_phase phase);
    //   super.start_of_simulation_phase(phase);
    //   uvm_test_top.print_topology(uvm_default_tree_printer);
    // endfunction
  
    virtual function void build_phase(uvm_phase phase);
      super.build_phase(phase);
      e0 = env::type_id::create("e0", this);
      if (!uvm_config_db#(virtual reg_if)::get(this, "", "reg_vif", vif))
        `uvm_fatal("TEST", "Did not get vif")
  
        uvm_config_db#(virtual reg_if)::set(this, "e0.a0.*", "reg_vif", vif);
    endfunction
  
    virtual task run_phase(uvm_phase phase);
      gen_item_seq seq = gen_item_seq::type_id::create("seq");
      phase.raise_objection(this);
      apply_reset();
  
      seq.randomize() with {num inside {[20:30]}; };
      seq.start(e0.a0.s0);
      #200;
      phase.drop_objection(this);
    endtask
  
    virtual task apply_reset();
      vif.rstn <= 0;
      repeat(5) @ (posedge vif.clk);
      vif.rstn <= 1;
      repeat(10) @ (posedge vif.clk);
    endtask
endclass